library IEEE;
use IEEE.std_logic_1164.all;

entity ShiftRegisterDemo is
    port (sw : in std_logic_vector)